`timescale 1ns / 1ps

module ROM (
    input logic [31:0] addr,

    output logic [31:0] data
);

    logic [31:0] rom[0:61];

    assign data = rom[addr[31:2]];      //32bit 단위 --> 4B단위로 주소 처리: 하위 2bit 없애면 4B단위 처리 가능
    
//////////////////////////////////TEST용
    initial begin
        //rom[x] = 32'b func7 _ rs2 _ rs1 _ func3 _ rd _ op
        rom[0] = 32'b0000000_00001_00010_000_00100_0110011;    //add x4, x2, x1 O
        rom[1] = 32'b0100000_00001_00010_000_00101_0110011;    //sub x5, x2, x1 O
        rom[2] = 32'b0000000_00001_00100_001_00110_0110011;    //sll x6, x4, x1 O
        rom[3] = 32'b0000000_00011_00101_101_00111_0110011;    //srl x7, x5, x3 O
        rom[4] = 32'b0100000_00010_01111_101_01000_0110011;    //sra x8, x15, x2
        rom[5] = 32'b0000000_01000_00111_010_01001_0110011;    //slt x9, x7, x8
        rom[6] = 32'b0000000_01110_01111_011_01010_0110011;    //sltu x10, x13, x12
        rom[7] = 32'b0000000_00001_00100_100_01011_0110011;    //xor x11, x4, x1
        rom[8] = 32'b0000000_00011_00010_110_01100_0110011;    //or x12, x2, x3
        rom[9] = 32'b0000000_00111_00101_111_01101_0110011;    //and x13, x5, x7
    end
//////////////////////////////////

endmodule
